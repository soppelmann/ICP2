//------------------------------------------------------------------------------
// clock_if interface
//
// This interface provides a clock output signal.
// 
//------------------------------------------------------------------------------
interface clock_if ();
    // clock output signal.
    logic clock;
endinterface : clock_if

